`include "mux16to1.v"
module rightshifter(A, S, Y);
   input [15:0] A;  // The value to be shifted.
   input [3:0] S;  // The amount to shift.
   output [15:0] Y;  // The shifted result.

   mux16to1 mux0(Y[0], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], S[3], S[2], S[1], S[0]);
   mux16to1 mux1(Y[1], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], S[3], S[2], S[1], S[0]);
   mux16to1 mux2(Y[2], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], S[3], S[2], S[1], S[0]);
   mux16to1 mux3(Y[3], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2],  S[3], S[2], S[1], S[0]);
   mux16to1 mux4(Y[4], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3],  S[3], S[2], S[1], S[0]);
   mux16to1 mux5(Y[5], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], S[3], S[2], S[1], S[0]);
   mux16to1 mux6(Y[6], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], S[3], S[2], S[1], S[0]);
   mux16to1 mux7(Y[7], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], S[3], S[2], S[1], S[0]);
   mux16to1 mux8(Y[8], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], S[3], S[2], S[1], S[0]);
   mux16to1 mux9(Y[9], A[9], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], S[3], S[2], S[1], S[0]);
   mux16to1 mux10(Y[10], A[10], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], S[3], S[2], S[1], S[0]);
   mux16to1 mux11(Y[11], A[11], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], S[3], S[2], S[1], S[0]);
   mux16to1 mux12(Y[12], A[12], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], S[3], S[2], S[1], S[0]);
   mux16to1 mux13(Y[13], A[13], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], S[3], S[2], S[1], S[0]);
   mux16to1 mux14(Y[14], A[14], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], S[3], S[2], S[1], S[0]);
   mux16to1 mux15(Y[15], A[15], A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], S[3], S[2], S[1], S[0]);
endmodule

module leftshifter(A, S, Y);
   input [15:0] A;  // The value to be shifted.
   input [3:0] S;  // The amount to shift.
   output [15:0] Y;  // The shifted result.

   mux16to1 mux0(Y[0], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], S[3], S[2], S[1], S[0]);
   mux16to1 mux1(Y[1], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], S[3], S[2], S[1], S[0]);
   mux16to1 mux2(Y[2], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], S[3], S[2], S[1], S[0]);
   mux16to1 mux3(Y[3], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4],  S[3], S[2], S[1], S[0]);
   mux16to1 mux4(Y[4], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5],  S[3], S[2], S[1], S[0]);
   mux16to1 mux5(Y[5], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], S[3], S[2], S[1], S[0]);
   mux16to1 mux6(Y[6], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], S[3], S[2], S[1], S[0]);
   mux16to1 mux7(Y[7], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], S[3], S[2], S[1], S[0]);
   mux16to1 mux8(Y[8], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], A[9], S[3], S[2], S[1], S[0]);
   mux16to1 mux9(Y[9], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], A[10], S[3], S[2], S[1], S[0]);
   mux16to1 mux10(Y[10], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], A[11], S[3], S[2], S[1], S[0]);
   mux16to1 mux11(Y[11], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], A[12], S[3], S[2], S[1], S[0]);
   mux16to1 mux12(Y[12], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], A[13], S[3], S[2], S[1], S[0]);
   mux16to1 mux13(Y[13], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], A[14], S[3], S[2], S[1], S[0]);
   mux16to1 mux14(Y[14], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], A[15], S[3], S[2], S[1], S[0]);
   mux16to1 mux15(Y[15], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], S[3], S[2], S[1], S[0]);
endmodule